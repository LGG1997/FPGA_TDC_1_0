`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/24/2021 09:12:56 AM
// Design Name: 
// Module Name: _48_6_encoder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//priority encoder
module _48_6_encoder
	#(
	 	parameter INDEX = 0
	)
	( 
	  input clk,
	  input rst,  
      input en,
      input [47:0] din,
      output reg [5:0] dout,
      output reg [9:0] offset,
      output reg Yen,
	  output reg Ynem
    );

reg [5:0] tmp;
reg [47:0]tmp_din;

always @(posedge clk or posedge rst) begin
    if(rst == 1'b1) begin
        tmp_din <= 0;
    end
    else begin
        tmp_din <= din;
    end
end


always @(*) begin
        casez(tmp_din)
        {{47{1'b0}},{1{1'b?}}}        :  tmp <= 6'b000000;  //48'b0000_0000_0000_0000_0000_0000_0000_000?
        {{46{1'b0}},1'b1,{1{1'b?}}}   :  tmp <= 6'b000001;  //48'b0000_0000_0000_0000_0000_0000_0000_001?
        {{45{1'b0}},1'b1,{2{1'b?}}}   :  tmp <= 6'b000010;  //48'b0000_0000_0000_0000_0000_0000_0000_01??
        {{44{1'b0}},1'b1,{3{1'b?}}}   :  tmp <= 6'b000011;  //48'b0000_0000_0000_0000_0000_0000_0000_1???
        {{43{1'b0}},1'b1,{4{1'b?}}}   :  tmp <= 6'b000100;  //48'b0000_0000_0000_0000_0000_0000_0001_????
        {{42{1'b0}},1'b1,{5{1'b?}}}   :  tmp <= 6'b000101;  //48'b0000_0000_0000_0000_0000_0000_001?_????
        {{41{1'b0}},1'b1,{6{1'b?}}}   :  tmp <= 6'b000110;  //48'b0000_0000_0000_0000_0000_0000_01??_????
        {{40{1'b0}},1'b1,{7{1'b?}}}   :  tmp <= 6'b000111;  //48'b0000_0000_0000_0000_0000_0000_1???_????
        {{39{1'b0}},1'b1,{8{1'b?}}}   :  tmp <= 6'b001000;  //48'b0000_0000_0000_0000_0000_0001_????_????
        {{38{1'b0}},1'b1,{9{11'b?}}}  :  tmp <= 6'b001001;  //48'b0000_0000_0000_0000_0000_001?_????_????
        {{37{1'b0}},1'b1,{10{1'b?}}}  :  tmp <= 6'b001010;  //48'b0000_0000_0000_0000_0000_01??_????_????
        {{36{1'b0}},1'b1,{11{1'b?}}}  :  tmp <= 6'b001011;  //48'b0000_0000_0000_0000_0000_1???_????_????
        {{35{1'b0}},1'b1,{12{1'b?}}}  :  tmp <= 6'b001100;  //48'b0000_0000_0000_0000_0001_????_????_????
        {{34{1'b0}},1'b1,{13{1'b?}}}  :  tmp <= 6'b001101;  //48'b0000_0000_0000_0000_001?_????_????_????
        {{33{1'b0}},1'b1,{15{1'b?}}}  :  tmp <= 6'b001110;  //48'b0000_0000_0000_0000_01??_????_????_????
        {{32{1'b0}},1'b1,{15{1'b?}}}  :  tmp <= 6'b001111;  //48'b0000_0000_0000_0000_1???_????_????_????
        
        {{31{1'b0}},1'b1,{16{1'b?}}}  :  tmp <= 6'b010000;  
        {{30{1'b0}},1'b1,{17{1'b?}}}  :  tmp <= 6'b010001;  
        {{29{1'b0}},1'b1,{18{1'b?}}}  :  tmp <= 6'b010010;  
        {{28{1'b0}},1'b1,{19{1'b?}}}  :  tmp <= 6'b010011;  
        {{27{1'b0}},1'b1,{20{1'b?}}}  :  tmp <= 6'b010100;  
        {{26{1'b0}},1'b1,{21{1'b?}}}  :  tmp <= 6'b010101;  
        {{25{1'b0}},1'b1,{22{1'b?}}}  :  tmp <= 6'b010110;  
        {{24{1'b0}},1'b1,{23{1'b?}}}  :  tmp <= 6'b010111;  
        {{23{1'b0}},1'b1,{24{1'b?}}}  :  tmp <= 6'b011000;  
        {{22{1'b0}},1'b1,{25{1'b?}}}  :  tmp <= 6'b011001;  
        {{21{1'b0}},1'b1,{26{1'b?}}}  :  tmp <= 6'b011010;  
        {{20{1'b0}},1'b1,{27{1'b?}}}  :  tmp <= 6'b011011; 
        {{19{1'b0}},1'b1,{28{1'b?}}}  :  tmp <= 6'b011100; 
        {{18{1'b0}},1'b1,{29{1'b?}}}  :  tmp <= 6'b011101;  
        {{17{1'b0}},1'b1,{30{1'b?}}}  :  tmp <= 6'b011110;  
        {{16{1'b0}},1'b1,{31{1'b?}}}  :  tmp <= 6'b011111; 
        
        {{15{1'b0}},1'b1,{32{1'b?}}}  :  tmp <= 6'b100000;  
        {{14{1'b0}},1'b1,{33{1'b?}}}  :  tmp <= 6'b100001;  
        {{13{1'b0}},1'b1,{34{1'b?}}}  :  tmp <= 6'b100010;  
        {{12{1'b0}},1'b1,{35{1'b?}}}  :  tmp <= 6'b100011;  
        {{11{1'b0}},1'b1,{36{1'b?}}}  :  tmp <= 6'b100100;  
        {{10{1'b0}},1'b1,{37{1'b?}}}  :  tmp <= 6'b100101;  
        {{9{1'b0}},1'b1,{38{1'b?}}}   :  tmp <= 6'b100110;  
        {{8{1'b0}},1'b1,{39{1'b?}}}   :  tmp <= 6'b100111;  
        {{7{1'b0}},1'b1,{40{1'b?}}}   :  tmp <= 6'b101000;  
        {{6{1'b0}},1'b1,{41{1'b?}}}   :  tmp <= 6'b101001;  
        {{5{1'b0}},1'b1,{42{1'b?}}}   :  tmp <= 6'b101010;  
        {{4{1'b0}},1'b1,{43{1'b?}}}   :  tmp <= 6'b101011; 
        {{3{1'b0}},1'b1,{44{1'b?}}}   :  tmp <= 6'b101100; 
        {{2{1'b0}},1'b1,{45{1'b?}}}   :  tmp <= 6'b101101;  
        {{1{1'b0}},1'b1,{46{1'b?}}}   :  tmp <= 6'b101110;  
        {{0{1'b0}},1'b1,{47{1'b?}}}   :  tmp <= 6'b101111; 
        default:
            tmp <= 6'b000000;
        endcase
   
end

always @(posedge clk or posedge rst) 
begin
	if(rst == 1) begin
		dout <= 0;
		Ynem <= 0;			
		Yen <=  0;
		offset <= 0;
	end
	else begin
		dout <= tmp;
		Ynem <= (tmp_din != {48{1'b0}}) ? 1'b1 : 1'b0;			
		Yen <=  (tmp_din == {48{1'b0}})? 1'b1 : 1'b0;
		offset <= (tmp_din != {48{1'b0}}) ? INDEX*48 : 10'b00_0000_0000;
	end
end

endmodule
